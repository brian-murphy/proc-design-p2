`ifndef _pc_apparatus_vh_
`define _pc_apparatus_vh_

`define PCSEL_PCPLUSFOUR 2'b00
`define PCSEL_PCOFFSET 2'b01
`define PCSEL_REGOFFSET 2'b10

`endif
