`ifndef _ui_controller_vh_
`define _ui_controller_vh_

`define UI_KEY 2'b00
`define UI_SW 2'b01
`define UI_LEDR 2'b10
`define UI_HEX 2'b11

`endif