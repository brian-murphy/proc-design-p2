`ifndef _alu_vh_
`define _alu_vh_

`define ADD 5'd0
`define SUB 5'd1
`define AND 5'd2
`define OR 5'd3
`define XOR 5'd4
`define NAND 5'd5
`define NOR 5'd6
`define XNOR 5'd7
`define MVHI 5'd8
`define F 5'd9
`define EQ 5'd10
`define LT 5'd11
`define LTE 5'd12
`define T 5'd13
`define NE 5'd14
`define GTE 5'd15
`define GT 5'd16

`define WORD_SIZE 32
`define FUNC_BITS 5

// `define M (`N << 2)
`endif
