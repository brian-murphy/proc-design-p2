`ifndef _io_controller_vh_
`define _io_controller_vh_

`define IO_LOAD 1'b0
`define IO_STORE 1'b1

`endif
