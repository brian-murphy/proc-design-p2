`ifndef _ui_controller_vh_
`define _ui_controller_vh_

`define KEY 2'b00
`define SW 2'b01
`define LEDR 2'b10
`define HEX 2'b11

`endif