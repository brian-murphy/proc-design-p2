`ifndef _alu_vh_
`define _alu_vh_

`define ADD 0
`define SUB 1
`define AND 2
`define OR 3
`define XOR 4
`define NAND 5
`define NOR 6
`define XNOR 7
`define MVHI 8
`define F 9
`define EQ 10
`define LT 11
`define LTE 12
`define T 13
`define NE 14
`define GTE 15
`define GT 16


// `define M (`N << 2)
`endif //_my_incl_vh_
